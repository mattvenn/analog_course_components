magic
tech sky130A
magscale 1 2
timestamp 1715860637
<< pwell >>
rect -739 -2582 739 2582
<< psubdiff >>
rect -703 2512 -607 2546
rect 607 2512 703 2546
rect -703 2450 -669 2512
rect 669 2450 703 2512
rect -703 -2512 -669 -2450
rect 669 -2512 703 -2450
rect -703 -2546 -607 -2512
rect 607 -2546 703 -2512
<< psubdiffcont >>
rect -607 2512 607 2546
rect -703 -2450 -669 2450
rect 669 -2450 703 2450
rect -607 -2546 607 -2512
<< xpolycontact >>
rect -573 1984 573 2416
rect -573 -2416 573 -1984
<< ppolyres >>
rect -573 -1984 573 1984
<< locali >>
rect -703 2512 -607 2546
rect 607 2512 703 2546
rect -703 2450 -669 2512
rect 669 2450 703 2512
rect -703 -2512 -669 -2450
rect 669 -2512 703 -2450
rect -703 -2546 -607 -2512
rect 607 -2546 703 -2512
<< viali >>
rect -557 2001 557 2398
rect -557 -2398 557 -2001
<< metal1 >>
rect -569 2398 569 2404
rect -569 2001 -557 2398
rect 557 2001 569 2398
rect -569 1995 569 2001
rect -569 -2001 569 -1995
rect -569 -2398 -557 -2001
rect 557 -2398 569 -2001
rect -569 -2404 569 -2398
<< properties >>
string FIXED_BBOX -686 -2529 686 2529
string gencell sky130_fd_pr__res_high_po_5p73
string library sky130
string parameters w 5.730 l 20.0 m 1 nx 1 wmin 5.730 lmin 0.50 rho 319.8 val 1.184k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 5.730 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
