** sch_path: /home/matt/work/asic-workshop/shuttle-2404/analog_course_components/xschem/res.sch
.subckt res r1_r0 r2_r0 r1_r1 r2_r1 subs
*.PININFO r1_r0:B r2_r0:B r1_r1:B r2_r1:B subs:B
XR1 r1_r1 r1_r0 subs sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR2 r2_r1 r2_r0 subs sky130_fd_pr__res_high_po_5p73 L=20 mult=1 m=1
.ends
.end
